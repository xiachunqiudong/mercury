package mercury_pkg;

  typedef struct packed {
    logic [4:0] lsrc1;
    logic [4:0] lsrc2;
    logic [4:0] ldst;
  } uop_info_t;

endpackage