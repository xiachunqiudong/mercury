module exu_decoder(
  input  logic [31:0] inst,
  output logic [4:0]  lsrc1,
  output logic [4:0]  lsrc2,
  output logic [4:0]  ldst
);



endmodule